library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
 
entity Modo is
    port (
        clk  : in std_logic;
        en   : in std_logic;
		  state: in std_logic_vector(1 downto 0);
        addr : in std_logic_vector(9 downto 0);
        data : out std_logic_vector(47 to 66)
    );
end modo;
 
architecture behavioral of modo is
    type memoria_rom is array (21 to 40) of std_logic_vector (47 to 66);
    signal Anim: memoria_rom;
	 signal ROM1 : memoria_rom := (
	 "11111111111111111111",
	 "10000000000000000001",
	 "10000111111111100001",
	 "10000111111111100001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10000111111111100001",
	 "10000111111111100001",
	 "10000000000000000001",
	 "11111111111111111111"
	 );
	signal ROM2 : memoria_rom := (
	 "11111111111111111111",
	 "10000000000000000001",
	 "10000000111100000001",
	 "10000001100110000001",
	 "10000011000011000001",
	 "10000011000011000001",
	 "10000110000001100001",
	 "10000110000001100001",
	 "10001100000000110001",
	 "10001100000000110001",
	 "10011000000000011001",
	 "10011111111111111001",
	 "10011111111111111001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10000000000000000001",
	 "11111111111111111111"
	 );
	 signal ROM3 : memoria_rom := (
	 "11111111111111111111",
	 "10000000000000000001",
	 "10000110000001100001",
	 "10000110000001100001",
	 "10011011000011011001",
	 "10011011000011011001",
	 "10011001100110011001",
	 "10011001100110011001",
	 "10011000011000011001",
	 "10011000011000011001",
	 "10011000011000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10011000000000011001",
	 "10000000000000000001",
	 "11111111111111111111"
	 );
begin
	 anim <= ROM3 when state = "10" else
				ROM3 when state = "11" else
				ROM3 when state = "00" else
				ROM3 when state = "01" else
				anim;
    process (clk) begin
        if rising_edge(clk) then
            if (en = '1') then
                if(addr >=21 and addr <=40) then
						data <= anim(conv_integer(addr));
					 else data <= (others=>'0');
					 end if;
            end if;
        end if;
    end process;
end behavioral;