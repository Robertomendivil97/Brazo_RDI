library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
 
entity claw_anim is
    port (
        clk  : in std_logic;
        en   : in std_logic;
		  state: in std_logic_vector(1 downto 0);
        addr : in std_logic_vector(9 downto 0);
        data : out std_logic_vector(401 to 592)
    );
end claw_anim;
 
architecture behavioral of claw_anim is
    type memoria_rom is array (287 to 438) of std_logic_vector (401 to 592);
    signal Anim: memoria_rom;
	 signal ROM1 : memoria_rom := (
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
	 );
	 signal ROM2 : memoria_rom := (
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
	 );
	 signal ROM3 : memoria_rom := (
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	 "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
	 );
begin
	 anim <= ROM1 when state = "00" else
				ROM2 when state = "01" else
				ROM3 when state = "10" else
				anim;
    process (clk) begin
        if rising_edge(clk) then
            if (en = '1') then
                if(addr >=287 and addr <=438) then
						data <= anim(conv_integer(addr));
					 else data <= (others=>'0');
					 end if;
            end if;
        end if;
    end process;
end behavioral;