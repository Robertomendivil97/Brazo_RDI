library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
 
entity motor1_estatus is
    port (
        clk  : in std_logic;
        en   : in std_logic;
		  state: in std_logic_vector(1 downto 0);
        addr : in std_logic_vector(9 downto 0);
        data : out std_logic_vector(47 to 86)
    );
end motor1_estatus;
 
architecture behavioral of motor1_estatus is
    type memoria_rom is array (43 to 102) of std_logic_vector (47 to 86);
    signal Anim: memoria_rom;
	 
	 signal ROM1 : memoria_rom := (
	 "1111111111111111111111111111111111111111",
	 "1000000000000000000000000000000000000001",
	 "1000011000000110000000000011111100000001",
	 "1000011000000110000000000111111100000001",
	 "1001101100001101100000001111111100000001",
	 "1001101100001101100000011111111100000001",
	 "1001100110011001100000000001111100000001",
	 "1001100110011001100000000001111100000001",
	 "1001100001100001100000000001111100000001",
	 "1001100001100001100000000001111100000001",
	 "1001100001100001100000000001111100000001",
	 "1001100000000001100000000001111100000001",
	 "1001100000000001100000000001111100000001",
	 "1001100000000001100000000001111100000001",
	 "1001100000000001100000000001111100000001",
	 "1001100000000001100000000001111100000001",
	 "1001100000000001100000111111111111111001",
	 "1001100000000001100000111111111111111001",
	 "1000000000000000000000000000000000000001",
	 "1111111111111111111111111111111111111111",
	 "1111111111111111111111111111111111111111",
	 "1000000000000000000000000000000000000001",
	 "1000011000000110000000000001111000000001",
	 "1000011000000110000000000011111100000001",
	 "1001101100001101100000000111001110000001",
	 "1001101100001101100000001110000111000001",
	 "1001100110011001100000011100000011100001",
	 "1001100110011001100000111000000001110001",
	 "1001100001100001100000000000000000111001",
	 "1001100001100001100000000000000000111001",
	 "1001100001100001100000000000000011100001",
	 "1001100000000001100000000000001110000001",
	 "1001100000000001100000000000111000000001",
	 "1001100000000001100000000011100000000001",
	 "1001100000000001100000001110000000000001",
	 "1001100000000001100000111000000000000001",
	 "1001100000000001100000111111111111111001",
	 "1001100000000001100000111111111111111001",
	 "1000000000000000000000000000000000000001",
	 "1111111111111111111111111111111111111111",
	 "1111111111111111111111111111111111111111",
	 "1000000000000000000000000000000000000001",
	 "1000011000000110000000111111111111000001",
	 "1000011000000110000000111111111111000001",
	 "1001101100001101100000111111111111000001",
	 "1001101100001101100000111111111111000001",
	 "1001100110011001100000000000011111111001",
	 "1001100110011001100000000000011111111001",
	 "1001100001100001100000111111111111000001",
	 "1001100001100001100000111111111111000001",
	 "1001100001100001100000111111111111000001",
	 "1001100000000001100000111111111111000001",
	 "1001100000000001100000000000011111111001",
	 "1001100000000001100000000000011111111001",
	 "1001100000000001100000111111111111000001",
	 "1001100000000001100000111111111111000001",
	 "1001100000000001100000111111111111000001",
	 "1001100000000001100000111111111111000001",
	 "1000000000000000000000000000000000000001",
	 "1111111111111111111111111111111111111111"
	 );
begin
	 anim <= ROM1;
    process (clk) begin
        if rising_edge(clk) then
            if (en = '1') then
                if(addr >=43 and addr <=102) then
						data <= anim(conv_integer(addr));
					 else data <= (others=>'0');
					 end if;
            end if;
        end if;
    end process;
end behavioral;
